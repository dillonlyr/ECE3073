
module NIOSII_WEEK2 (
	clk_clk,
	led_export,
	reset_reset_n,
	gpio_export);	

	input		clk_clk;
	output	[7:0]	led_export;
	input		reset_reset_n;
	output		gpio_export;
endmodule
